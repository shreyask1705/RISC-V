module testbench_riscv



endmodule